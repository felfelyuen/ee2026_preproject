`timescale 1ns / 1ps

//////////////////////////////////////////////////////////////////////////////////
//
//  FILL IN THE FOLLOWING INFORMATION:
//  STUDENT A NAME: 
//  STUDENT B NAME:
//  STUDENT C NAME: 
//  STUDENT D NAME:  
//
//////////////////////////////////////////////////////////////////////////////////

module Top_Student (
    input CLK,
    input CTRLbtn, 
    input UPbtn,
    input DOWNbtn,
    output [7:0] Jx
    );
        task_B task2 (CLK, CTRLbtn, UPbtn, DOWNbtn);
endmodule
